/////////////////////////////////////////////////////////////////////////
//                                                                     //
//   Modulename :  cpu.sv                                              //
//                                                                     //
//  Description :  Top-level module of the verisimple processor;       //
//                 This instantiates and connects the 5 stages of the  //
//                 Verisimple pipeline together.                       //
//                                                                     //
/////////////////////////////////////////////////////////////////////////

`include "sys_defs.svh"

module cpu (
    input clock, // System clock
    input reset, // System reset

    input MEM_TAG   mem2proc_transaction_tag, // Memory tag for current transaction
    input MEM_BLOCK mem2proc_data,            // Data coming back from memory
    input MEM_TAG   mem2proc_data_tag,        // Tag for which transaction data is for

    output MEM_COMMAND proc2mem_command, // Command sent to memory
    output ADDR        proc2mem_addr,    // Address sent to memory
    output MEM_BLOCK   proc2mem_data,    // Data sent to memory
    output MEM_SIZE    proc2mem_size,    // Data size sent to memory

    // Note: these are assigned at the very bottom of the module
    output COMMIT_PACKET [`N-1:0] committed_insts,

    // Debug outputs: these signals are solely used for debugging in testbenches
    // Do not change for project 3
    // You should definitely change these for project 4
    output ADDR  if_NPC_dbg,
    output DATA  if_inst_dbg,
    output logic if_valid_dbg,
    output ADDR  if_id_NPC_dbg,
    output DATA  if_id_inst_dbg,
    output logic if_id_valid_dbg,
    output ADDR  id_ex_NPC_dbg,
    output DATA  id_ex_inst_dbg,
    output logic id_ex_valid_dbg,
    output ADDR  ex_mem_NPC_dbg,
    output DATA  ex_mem_inst_dbg,
    output logic ex_mem_valid_dbg,
    output ADDR  mem_wb_NPC_dbg,
    output DATA  mem_wb_inst_dbg,
    output logic mem_wb_valid_dbg
);

    //////////////////////////////////////////////////
    //                                              //
    //                Pipeline Wires                //
    //                                              //
    //////////////////////////////////////////////////

    // Pipeline register enables
    logic if_id_enable, id_ex_enable, ex_mem_enable, mem_wb_enable;

    // Outputs from IF-Stage and IF/ID Pipeline Register
    ADDR Imem_addr;
    IF_ID_PACKET if_packet, if_id_reg;

    // Outputs from ID stage and ID/EX Pipeline Register
    ID_EX_PACKET id_packet, id_ex_reg;

    // Outputs from EX-Stage and EX/MEM Pipeline Register
    EX_MEM_PACKET ex_packet, ex_mem_reg;

    // Outputs from MEM-Stage and MEM/WB Pipeline Register
    MEM_WB_PACKET mem_packet, mem_wb_reg;

    // Outputs from MEM-Stage to memory
    ADDR        Dmem_addr;
    MEM_BLOCK   Dmem_store_data;
    MEM_COMMAND Dmem_command;
    MEM_SIZE    Dmem_size;

    // Outputs from WB-Stage (These loop back to the register file in ID)
    COMMIT_PACKET wb_packet;

    // forwarding unit
    logic [1:0] forward_a, forward_b;

    // control unit
    logic flush;

    // stall
    logic stall;

    //////////////////////////////////////////////////
    //                                              //
    //              structural hazard               //
    //                                              //
    //////////////////////////////////////////////////

    logic hazard_rs1;
    logic hazard_rs2;
    logic hazard_branch;
    logic hazard_store;

    assign hazard_rs1 = (id_packet.opa_select == OPA_IS_RS1) & (id_ex_reg.dest_reg_idx == id_packet.inst.r.rs1);
    assign hazard_rs2 = (id_packet.opb_select == OPB_IS_RS2) & (id_ex_reg.dest_reg_idx == id_packet.inst.r.rs2);
    assign hazard_branch = id_packet.cond_branch
                    & ((id_ex_reg.dest_reg_idx == id_packet.inst.r.rs1)
                    |  (id_ex_reg.dest_reg_idx == id_packet.inst.r.rs2));
    assign hazard_store = id_packet.wr_mem & (id_ex_reg.dest_reg_idx == id_packet.inst.s.rs2);
    assign stall = id_ex_reg.valid & id_packet.valid & id_ex_reg.rd_mem & (id_ex_reg.dest_reg_idx != `ZERO_REG) & (hazard_branch | hazard_rs1 | hazard_rs2 | hazard_store);

    //////////////////////////////////////////////////
    //                                              //
    //                forward                       //
    //                                              //
    //////////////////////////////////////////////////

    always_comb begin
        forward_a = 2'b00;
        forward_b = 2'b00;

        if (ex_mem_reg.valid & !ex_mem_reg.rd_mem & (ex_mem_reg.dest_reg_idx != `ZERO_REG) & (ex_mem_reg.dest_reg_idx == id_ex_reg.inst.r.rs1)) begin
            forward_a = 2'b01;
        end else if (mem_wb_reg.valid & (mem_wb_reg.dest_reg_idx != `ZERO_REG) & (mem_wb_reg.dest_reg_idx == id_ex_reg.inst.r.rs1)) begin
            forward_a = 2'b10;
        end

        if (ex_mem_reg.valid & !ex_mem_reg.rd_mem & (ex_mem_reg.dest_reg_idx != `ZERO_REG) & (ex_mem_reg.dest_reg_idx == id_ex_reg.inst.r.rs2)) begin
            forward_b = 2'b01;
        end else if (mem_wb_reg.valid & (mem_wb_reg.dest_reg_idx != `ZERO_REG) & (mem_wb_reg.dest_reg_idx == id_ex_reg.inst.r.rs2)) begin
            forward_b = 2'b10;
        end
    end

    //////////////////////////////////////////////////
    //                                              //
    //                contral hazard                //
    //                                              //
    //////////////////////////////////////////////////

    // assign flush = ex_mem_reg.valid & ex_mem_reg.take_branch;
    assign flush = ex_mem_reg.take_branch;

    //////////////////////////////////////////////////
    //                                              //
    //                Memory Outputs                //
    //                                              //
    //////////////////////////////////////////////////

    // these signals go to and from the processor and memory
    // we give precedence to the mem stage over instruction fetch
    // note that there is no latency in project 3
    // but there will be a 100ns latency in project 4

    always_comb begin
        if (Dmem_command != MEM_NONE) begin  // read or write DATA from memory
            proc2mem_command = Dmem_command;
            proc2mem_size    = Dmem_size;   // size is never DOUBLE in project 3
            proc2mem_addr    = Dmem_addr;
        end else begin                      // read an INSTRUCTION from memory
            proc2mem_command = MEM_LOAD;
            proc2mem_addr    = Imem_addr;
            proc2mem_size    = DOUBLE;      // instructions load a full memory line (64 bits)
        end
        proc2mem_data = Dmem_store_data;
    end

    //////////////////////////////////////////////////
    //                                              //
    //                  Valid Bit                   //
    //                                              //
    //////////////////////////////////////////////////

    // This state controls the stall signal that artificially forces IF
    // to stall until the previous instruction has completed.
    // For project 3, start by assigning if_valid to always be 1

    logic if_valid, start_valid_on_reset, wb_valid;


    always_ff @(posedge clock) begin
        // Start valid on reset. Other stages (ID,EX,MEM,WB) start as invalid
        // Using a separate always_ff is necessary since if_valid is combinational
        // Assigning if_valid = reset doesn't work as you'd hope :/
        start_valid_on_reset <= reset;
    end

    // valid bit will cycle through the pipeline and come back from the wb stage
    // assign if_valid = start_valid_on_reset | wb_valid;
    assign if_valid = (~stall) & (~(ex_mem_reg.rd_mem | ex_mem_reg.wr_mem));

    //////////////////////////////////////////////////
    //                                              //
    //                  IF-Stage                    //
    //                                              //
    //////////////////////////////////////////////////

    stage_if stage_if_0 (
        // Inputs
        .clock (clock),
        .reset (reset),
        .if_valid      (if_valid),
        .take_branch   (ex_mem_reg.take_branch),
        .branch_target (ex_mem_reg.alu_result),
        .Imem_data     (mem2proc_data),

        // Outputs
        .if_packet (if_packet),
        .Imem_addr (Imem_addr)
    );

    // debug outputs
    assign if_NPC_dbg   = if_packet.NPC;
    assign if_inst_dbg  = if_packet.inst;
    assign if_valid_dbg = if_packet.valid;

    //////////////////////////////////////////////////
    //                                              //
    //            IF/ID Pipeline Register           //
    //                                              //
    //////////////////////////////////////////////////

    assign if_id_enable = ~stall;

    always_ff @(posedge clock) begin
        if (reset) begin
            if_id_reg.inst  <= `NOP;
            if_id_reg.valid <= `FALSE;
            if_id_reg.NPC   <= 0;
            if_id_reg.PC    <= 0;
        end else if(flush) begin
            if_id_reg.inst  <= `NOP;
            if_id_reg.valid <= `FALSE;
        end else if (if_id_enable) begin
            if_id_reg <= if_packet;
        end
    end

    // debug outputs
    assign if_id_NPC_dbg   = if_id_reg.NPC;
    assign if_id_inst_dbg  = if_id_reg.inst;
    assign if_id_valid_dbg = if_id_reg.valid;

    //////////////////////////////////////////////////
    //                                              //
    //                  ID-Stage                    //
    //                                              //
    //////////////////////////////////////////////////

    stage_id stage_id_0 (
        // Inputs
        .clock (clock),
        .reset (reset),
        .if_id_reg       (if_id_reg),
        .wb_regfile_en   (wb_packet.valid),
        .wb_regfile_idx  (wb_packet.reg_idx),
        .wb_regfile_data (wb_packet.data),

        // Output
        .id_packet (id_packet)
    );

    //////////////////////////////////////////////////
    //                                              //
    //            ID/EX Pipeline Register           //
    //                                              //
    //////////////////////////////////////////////////

    assign id_ex_enable = 1'b1;

    always_ff @(posedge clock) begin
        if (reset | flush) begin
            id_ex_reg <= '{
                `NOP, // we can't simply assign 0 because NOP is non-zero
                32'b0, // PC
                32'b0, // NPC
                32'b0, // rs1 select
                32'b0, // rs2 select
                OPA_IS_RS1,
                OPB_IS_RS2,
                `ZERO_REG,
                ALU_ADD,
                1'b0, // mult
                1'b0, // rd_mem
                1'b0, // wr_mem
                1'b0, // cond
                1'b0, // uncond
                1'b0, // halt
                1'b0, // illegal
                1'b0, // csr_op
                1'b0  // valid
            };
        end else if (id_ex_enable) begin
            if(stall) begin
                id_ex_reg <= '{
                    `NOP, // we can't simply assign 0 because NOP is non-zero
                    32'b0, // PC
                    32'b0, // NPC
                    32'b0, // rs1 select
                    32'b0, // rs2 select
                    OPA_IS_RS1,
                    OPB_IS_RS2,
                    `ZERO_REG,
                    ALU_ADD,
                    1'b0, // mult
                    1'b0, // rd_mem
                    1'b0, // wr_mem
                    1'b0, // cond
                    1'b0, // uncond
                    1'b0, // halt
                    1'b0, // illegal
                    1'b0, // csr_op
                    1'b0  // valid
                };
            end else begin
                id_ex_reg <= id_packet;
            end
        end
    end

    // debug outputs
    assign id_ex_NPC_dbg   = id_ex_reg.NPC;
    assign id_ex_inst_dbg  = id_ex_reg.inst;
    assign id_ex_valid_dbg = id_ex_reg.valid;

    //////////////////////////////////////////////////
    //                                              //
    //                  EX-Stage                    //
    //                                              //
    //////////////////////////////////////////////////
    
    logic [31:0] fwd_rs1, fwd_rs2;

    always_comb begin
        fwd_rs1 = id_ex_reg.rs1_value;
        fwd_rs2 = id_ex_reg.rs2_value;

        case (forward_a)
            2'b01: fwd_rs1 = ex_mem_reg.alu_result;
            2'b10: fwd_rs1 = mem_wb_reg.result;
            default: begin
                //
            end
        endcase

        case (forward_b)
            2'b01: fwd_rs2 = ex_mem_reg.alu_result;
            2'b10: fwd_rs2 = mem_wb_reg.result;
            default: begin
                //
            end
        endcase
    end
    ID_EX_PACKET id_ex_reg_fwd;
    always_comb begin
        id_ex_reg_fwd         = id_ex_reg;
        id_ex_reg_fwd.rs1_value = fwd_rs1;
        id_ex_reg_fwd.rs2_value = fwd_rs2;
    end


    stage_ex stage_ex_0 (
        // Input
        .id_ex_reg (id_ex_reg_fwd),

        // Output
        .ex_packet (ex_packet)
    );

    //////////////////////////////////////////////////
    //                                              //
    //           EX/MEM Pipeline Register           //
    //                                              //
    //////////////////////////////////////////////////

    assign ex_mem_enable = 1'b1;

    always_ff @(posedge clock) begin
        if (reset | flush) begin
            ex_mem_inst_dbg <= `NOP; // debug output
            ex_mem_reg      <= 0;    // the defaults can all be zero!
        end else if (ex_mem_enable) begin
            ex_mem_inst_dbg <= id_ex_inst_dbg; // debug output, just forwarded from ID
            ex_mem_reg      <= ex_packet;
        end
    end

    // debug outputs
    assign ex_mem_NPC_dbg   = ex_mem_reg.NPC;
    assign ex_mem_valid_dbg = ex_mem_reg.valid;

    //////////////////////////////////////////////////
    //                                              //
    //                 MEM-Stage                    //
    //                                              //
    //////////////////////////////////////////////////

    stage_mem stage_mem_0 (
        // Inputs
        .ex_mem_reg     (ex_mem_reg),
        .Dmem_load_data (mem2proc_data),

        // Outputs
        .mem_packet      (mem_packet),
        .Dmem_command    (Dmem_command),
        .Dmem_size       (Dmem_size),
        .Dmem_addr       (Dmem_addr),
        .Dmem_store_data (Dmem_store_data)
    );

    //////////////////////////////////////////////////
    //                                              //
    //           MEM/WB Pipeline Register           //
    //                                              //
    //////////////////////////////////////////////////

    assign mem_wb_enable = 1'b1;

    always_ff @(posedge clock) begin
        if (reset) begin
            mem_wb_inst_dbg <= `NOP; // debug output
            mem_wb_reg      <= 0;    // the defaults can all be zero!
        end else if (mem_wb_enable) begin
            mem_wb_inst_dbg <= ex_mem_inst_dbg; // debug output, just forwarded from EX
            mem_wb_reg      <= mem_packet;
        end
    end

    // debug outputs
    assign mem_wb_NPC_dbg   = mem_wb_reg.NPC;
    assign mem_wb_valid_dbg = mem_wb_reg.valid;

    //////////////////////////////////////////////////
    //                                              //
    //                  WB-Stage                    //
    //                                              //
    //////////////////////////////////////////////////

    stage_wb stage_wb_0 (
        // Input
        .mem_wb_reg (mem_wb_reg), // doesn't use all of these

        // Output
        .wb_packet (wb_packet)
    );

    // This signal is solely used by if_valid for the initial stalling behavior
    always_ff @(posedge clock) begin
        if (reset) wb_valid <= 0;
        else       wb_valid <= mem_wb_reg.valid;
    end

    //////////////////////////////////////////////////
    //                                              //
    //               Pipeline Outputs               //
    //                                              //
    //////////////////////////////////////////////////

    // Output the committed instruction to the testbench for counting
    assign committed_insts[0] = wb_packet;

endmodule // pipeline